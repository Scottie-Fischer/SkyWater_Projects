magic
tech sky130A
timestamp 1647385306
<< nwell >>
rect -52 76 256 237
<< pwell >>
rect -52 -95 256 76
<< nmos >>
rect 0 0 15 42
rect 188 0 203 42
<< scnmos >>
rect 25 -49 61 -34
rect 142 -49 178 -34
<< pmos >>
rect 0 161 15 203
rect 188 161 203 203
<< ndiff >>
rect -29 29 0 42
rect -29 12 -25 29
rect -8 12 0 29
rect -29 0 0 12
rect 15 36 61 42
rect 15 19 38 36
rect 55 19 61 36
rect 15 0 61 19
rect 142 36 188 42
rect 142 19 148 36
rect 165 19 188 36
rect 25 -34 61 0
rect 142 0 188 19
rect 203 29 232 42
rect 203 12 211 29
rect 228 12 232 29
rect 203 0 232 12
rect 142 -34 178 0
rect 25 -58 61 -49
rect 25 -75 29 -58
rect 57 -75 61 -58
rect 25 -81 61 -75
rect 142 -58 178 -49
rect 142 -75 146 -58
rect 174 -75 178 -58
rect 142 -81 178 -75
<< pdiff >>
rect -27 192 0 203
rect -27 175 -23 192
rect -6 175 0 192
rect -27 161 0 175
rect 15 182 61 203
rect 15 165 38 182
rect 55 165 61 182
rect 15 161 61 165
rect 142 182 188 203
rect 142 165 148 182
rect 165 165 188 182
rect 142 161 188 165
rect 203 192 231 203
rect 203 175 210 192
rect 227 175 231 192
rect 203 161 231 175
<< ndiffc >>
rect -25 12 -8 29
rect 38 19 55 36
rect 148 19 165 36
rect 211 12 228 29
rect 29 -75 57 -58
rect 146 -75 174 -58
<< pdiffc >>
rect -23 175 -6 192
rect 38 165 55 182
rect 148 165 165 182
rect 210 175 227 192
<< poly >>
rect 0 203 15 216
rect 188 203 203 216
rect 0 72 15 161
rect 188 144 203 161
rect 40 136 203 144
rect 40 119 48 136
rect 65 129 203 136
rect 65 119 73 129
rect 40 111 73 119
rect 130 82 163 90
rect 130 72 138 82
rect 0 65 138 72
rect 155 65 163 82
rect 0 57 163 65
rect 0 42 15 57
rect 188 42 203 129
rect 0 -13 15 0
rect 82 6 121 14
rect 82 -17 90 6
rect 113 -17 121 6
rect 82 -34 121 -17
rect 188 -13 203 0
rect -52 -49 25 -34
rect 61 -49 142 -34
rect 178 -49 256 -34
<< polycont >>
rect 48 119 65 136
rect 138 65 155 82
rect 90 -17 113 6
<< locali >>
rect -52 227 256 237
rect -52 216 98 227
rect -25 213 98 216
rect -25 192 -6 213
rect 86 210 98 213
rect 115 216 256 227
rect 115 213 227 216
rect 115 210 124 213
rect 86 207 124 210
rect -25 175 -23 192
rect -25 167 -6 175
rect 38 182 61 196
rect 55 165 61 182
rect -52 144 -22 145
rect -52 125 -42 144
rect -25 125 -22 144
rect -52 124 -22 125
rect 38 144 61 165
rect 142 182 165 196
rect 142 165 148 182
rect 210 192 227 213
rect 210 167 227 175
rect 38 136 73 144
rect 38 119 48 136
rect 65 119 73 136
rect 38 111 73 119
rect -52 54 -43 71
rect -26 54 -22 71
rect -52 37 -22 54
rect -52 29 -8 37
rect -52 12 -25 29
rect -52 4 -8 12
rect 38 36 61 111
rect 142 90 165 165
rect 225 144 256 145
rect 225 125 228 144
rect 245 125 256 144
rect 225 124 256 125
rect 130 82 165 90
rect 130 65 138 82
rect 155 65 165 82
rect 130 57 165 65
rect 55 19 61 36
rect 38 11 61 19
rect 142 36 165 57
rect 225 54 229 71
rect 246 54 256 71
rect 225 37 256 54
rect 142 19 148 36
rect 82 7 121 14
rect 142 11 165 19
rect 211 29 256 37
rect 228 12 256 29
rect 82 -18 89 7
rect 114 -18 121 7
rect 211 4 256 12
rect 82 -25 121 -18
rect -2 -58 65 -56
rect -2 -75 -1 -58
rect 16 -75 29 -58
rect 57 -75 65 -58
rect -2 -77 65 -75
rect 138 -58 205 -56
rect 138 -75 146 -58
rect 174 -75 187 -58
rect 204 -75 205 -58
rect 138 -77 205 -75
<< viali >>
rect 98 210 115 227
rect -42 125 -25 144
rect -43 54 -26 71
rect 228 125 245 144
rect 229 54 246 71
rect 89 6 114 7
rect 89 -17 90 6
rect 90 -17 113 6
rect 113 -17 114 6
rect 89 -18 114 -17
rect -1 -75 16 -58
rect 187 -75 204 -58
<< metal1 >>
rect -52 144 -22 237
rect -52 125 -42 144
rect -25 125 -22 144
rect -52 71 -22 125
rect -52 54 -43 71
rect -26 54 -22 71
rect -52 -48 -22 54
rect -52 -74 -49 -48
rect -23 -74 -22 -48
rect -52 -95 -22 -74
rect -4 -58 19 237
rect 86 229 124 237
rect 86 202 92 229
rect 119 202 124 229
rect 86 199 124 202
rect 83 8 120 13
rect 83 -19 88 8
rect 115 -19 120 8
rect 83 -21 120 -19
rect -4 -75 -1 -58
rect 16 -75 19 -58
rect -4 -95 19 -75
rect 184 -58 207 237
rect 184 -75 187 -58
rect 204 -75 207 -58
rect 184 -95 207 -75
rect 225 144 256 237
rect 225 125 228 144
rect 245 125 256 144
rect 225 71 256 125
rect 225 54 229 71
rect 246 54 256 71
rect 225 -48 256 54
rect 225 -74 227 -48
rect 253 -74 256 -48
rect 225 -95 256 -74
<< via1 >>
rect -49 -74 -23 -48
rect 92 227 119 229
rect 92 210 98 227
rect 98 210 115 227
rect 115 210 119 227
rect 92 202 119 210
rect 88 7 115 8
rect 88 -18 89 7
rect 89 -18 114 7
rect 114 -18 115 7
rect 88 -19 115 -18
rect 227 -74 253 -48
<< metal2 >>
rect -52 229 256 237
rect -52 216 92 229
rect 86 202 92 216
rect 119 216 256 229
rect 119 202 124 216
rect 86 199 124 202
rect 85 8 118 11
rect 85 -19 88 8
rect 115 -19 118 8
rect 85 -20 118 -19
rect -52 -34 256 -20
rect -52 -74 -49 -48
rect -23 -74 227 -48
rect 253 -74 256 -48
rect -52 -77 256 -74
<< labels >>
rlabel polycont 48 119 65 136 1 q
rlabel polycont 138 65 155 82 1 qb
rlabel metal2 -52 -34 256 -20 1 wl
port 7 n
rlabel metal1 -4 -95 19 237 1 bl
port 1 n
rlabel metal1 184 -95 207 237 1 br
port 2 n
rlabel nwell -52 76 256 237 1 VPB
port 5 n
rlabel pwell -52 -95 256 76 1 VNB
port 6 n
rlabel metal2 -52 216 92 237 1 VPWR
port 4 n
rlabel metal1 -52 -95 -22 237 1 VGND
port 3 n
rlabel metal1 225 -95 256 237 1 VGND
<< end >>
